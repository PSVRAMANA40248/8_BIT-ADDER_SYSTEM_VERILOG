interface intf;
    logic [7:0] a, b;
    logic c;
    logic [7:0] sum;
    logic carry;
endinterface
